// ALU SIGNALS
