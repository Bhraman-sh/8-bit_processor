// INSTRUCTIONS OPCODE

`define MOV_A_B 8'h00
`define MOV_A_C 8'h01
`define MOV_A_D 8'h02

`define MOV_B_A 8'h03
`define MOV_B_C 8'h04
`define MOV_B_D 8'h05

`define MOV_C_B 8'h06
`define MOV_C_A 8'h07
`define MOV_C_D 8'h08

`define MOV_D_B 8'h09
`define MOV_D_C 8'h0a
`define MOV_D_A 8'h0b
