// CONTROLLER STATES

`define fetch         3'b000
`define decode        3'b001
`define execute       3'b010
`define store         3'b011
`define operand_fetch 3'b011
